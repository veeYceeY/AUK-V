library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;


entity code_mem is
    port(
            i_en : in std_logic;
            i_addr : in std_logic_vector(31 downto 0);
            o_data : out std_logic_vector(31 downto 0);
            o_valid: out std_logic
    );

end code_mem;

architecture behave of code_mem is
attribute rom_style : string;
type mem_type is array(1023 downto 0) of std_logic_vector(31 downto 0);
signal mem : mem_type;
attribute rom_style of mem : signal is "block";

begin
mem(6)<=x"07C00113";
mem(7)<=x"008000EF";
mem(8)<=x"0000006F";
mem(9)<=x"FD810113";
mem(10)<=x"02112223";
mem(11)<=x"02812023";
mem(12)<=x"02810413";
mem(13)<=x"07000793";
mem(14)<=x"FEF42423";
mem(15)<=x"07400793";
mem(16)<=x"FEF42223";
mem(17)<=x"07800793";
mem(18)<=x"FEF42023";
mem(19)<=x"FE842783";
mem(20)<=x"00500713";
mem(21)<=x"00E7A023";
mem(22)<=x"FE442783";
mem(23)<=x"00A00713";
mem(24)<=x"00E7A023";
mem(25)<=x"FE842783";
mem(26)<=x"0007A703";
mem(27)<=x"FE442783";
mem(28)<=x"0007A783";
mem(29)<=x"00F70733";
mem(30)<=x"FE042783";
mem(31)<=x"00E7A023";
mem(32)<=x"000017B7";
mem(33)<=x"00178793";
mem(34)<=x"FCF42E23";
mem(35)<=x"FDC42783";
mem(36)<=x"08600713";
mem(37)<=x"00E7A023";
mem(38)<=x"FE042A23";
mem(39)<=x"0100006F";
mem(40)<=x"FF442783";
mem(41)<=x"00178793";
mem(42)<=x"FEF42A23";
mem(43)<=x"FF442703";
mem(44)<=x"000317B7";
mem(45)<=x"D3F78793";
mem(46)<=x"FEE7D4E3";
mem(47)<=x"04500593";
mem(48)<=x"FDC42503";
mem(49)<=x"068000EF";
mem(50)<=x"FE042823";
mem(51)<=x"0100006F";
mem(52)<=x"FF042783";
mem(53)<=x"00178793";
mem(54)<=x"FEF42823";
mem(55)<=x"FF042703";
mem(56)<=x"000497B7";
mem(57)<=x"3DF78793";
mem(58)<=x"FEE7D4E3";
mem(59)<=x"07600593";
mem(60)<=x"FDC42503";
mem(61)<=x"038000EF";
mem(62)<=x"FE042623";
mem(63)<=x"0100006F";
mem(64)<=x"FEC42783";
mem(65)<=x"00178793";
mem(66)<=x"FEF42623";
mem(67)<=x"FEC42703";
mem(68)<=x"000317B7";
mem(69)<=x"D3F78793";
mem(70)<=x"FEE7D4E3";
mem(71)<=x"0E300593";
mem(72)<=x"FDC42503";
mem(73)<=x"008000EF";
mem(74)<=x"F71FF06F";
mem(75)<=x"FF010113";
mem(76)<=x"00812623";
mem(77)<=x"01010413";
mem(78)<=x"FEA42A23";
mem(79)<=x"FEB42823";
mem(80)<=x"FF442783";
mem(81)<=x"FF042703";
mem(82)<=x"00E7A023";
mem(83)<=x"00000013";
mem(84)<=x"00C12403";
mem(85)<=x"01010113";
mem(86)<=x"00008067";





--mem(0) <=x"03000413";
--mem(1) <=x"04000793";
--mem(2) <=x"FEF42623";
--mem(3) <=x"04400793";
--mem(4) <=x"FEF42423";
--mem(5) <=x"04800793";
--mem(6) <=x"FEF42223";
--mem(7) <=x"FE842783";
--mem(8) <=x"00A00713";
--mem(9) <=x"00E7A023";
--mem(10)<=x"FEC42783";
--mem(11)<=x"00400713";
--mem(12)<=x"00E7A023";
--mem(13)<=x"FEC42783";
--mem(14)<=x"0007A703";
--mem(15)<=x"FE842783";
--mem(16)<=x"0007A783";
--mem(17)<=x"00F70733";
--mem(18)<=x"FE442783";
--mem(19)<=x"00E7A023";
--mem(20)<=x"0000006F";

--working woith loops ---------
--mem(54)<=x"03000413";--
--mem(55)<=x"04000793";
--mem(56)<=x"FEF42023";
--mem(57)<=x"04400793";
--mem(58)<=x"FCF42E23";
--mem(59)<=x"04800793";
--mem(60)<=x"FCF42C23";
--mem(61)<=x"FE042783";
--mem(62)<=x"00500713";
--mem(63)<=x"00E7A023";
--mem(64)<=x"FDC42783";
--mem(65)<=x"00A00713";
--mem(66)<=x"00E7A023";
--mem(67)<=x"FE042783";
--mem(68)<=x"0007A703";
--mem(69)<=x"FDC42783";
--mem(70)<=x"0007A783";
--mem(71)<=x"00F70733";
--mem(72)<=x"FD842783";
--mem(73)<=x"00E7A023";
--mem(74)<=x"000017B7";
--mem(75)<=x"00178793";
--mem(76)<=x"FCF42A23";
--mem(77)<=x"FD442783";
--mem(78)<=x"08600713";
--mem(79)<=x"00E7A023";
--mem(80)<=x"FE042623";
--mem(81)<=x"FEC42703";
--mem(82)<=x"000317B7";
--mem(83)<=x"D3F78793";
--mem(84)<=x"00E7CA63";
--mem(85)<=x"FEC42783";
--mem(86)<=x"00178793";
--mem(87)<=x"FEF42623";
--mem(88)<=x"FE5FF06F";
--mem(89)<=x"FD442783";
--mem(90)<=x"04500713";
--mem(91)<=x"00E7A023";
--mem(92)<=x"FE042423";
--mem(93)<=x"FE842703";
--mem(94)<=x"000317B7";
--mem(95)<=x"D3F78793";
--mem(96)<=x"00E7CA63";
--mem(97)<=x"FE842783";
--mem(98)<=x"00178793";
--mem(99)<=x"FEF42423";
--mem(100)<=x"FE5FF06F";
--mem(101)<=x"FD442783";
--mem(102)<=x"07600713";
--mem(103)<=x"00E7A023";
--mem(104)<=x"FE042223";
--mem(105)<=x"FE442703";
--mem(106)<=x"000317B7";
--mem(107)<=x"D3F78793";
--mem(108)<=x"00E7CA63";
--mem(109)<=x"FE442783";
--mem(110)<=x"00178793";
--mem(111)<=x"FEF42223";
--mem(112)<=x"FE5FF06F";
--mem(113)<=x"FD442783";
--mem(114)<=x"0E300713";
--mem(115)<=x"00E7A023";
--mem(116)<=x"F71FF06F";


--     --        
     
-- mem(0) <= x"00044" & "00100" & "0110111";--LUI r1,#00044000h
-- mem(1) <= x"00032" & "00101" & "0110111";--LUI r2,#00032000h
-- mem(2) <= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R1,12
-- mem(3) <= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R2,12
-- mem(4) <= "0000000" & "00101" &"00100" &"000" & "00011" & "0110011";--ADD r3,r1,r2
-- mem(5) <= x"0000a" & "00001" & "0110111";--LUI r1,#00044000h
-- mem(6) <= x"00003" & "00010" & "0110111";--LUI r2,#00032000h
-- mem(7) <= "0000000" & "01100" &"00001" &"101" & "00001" & "0010011";--srlI R1,12
-- mem(8) <= "0000000" & "01100" &"00010" &"101" & "00010" & "0010011";--srlI R2,12
-- mem(9) <= x"0000f" & "00100" & "0110111";--LUI r4,0x0000a000
-- mem(10)<= x"00002" & "00101" & "0110111";--LUI r5,0x00004000
-- mem(11)<= x"00001" & "00110" & "0110111";--LUI r6,0x00001000
-- mem(12)<= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R4,12
-- mem(13)<= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R5,12
-- mem(14) <="0000000" & "01100" &"00110" &"101" & "00110" & "0010011";--srlI R6,12
-- mem(15) <= "0100000" & "00110" &"00100" &"000" & "00100" & "0110011";--sub r4,r4,r6
-- mem(16) <= "1111111" & "00100" &"00101" &"100" & "11101" & "1100011";--blt r4,r5,-1
-- mem(17) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(18) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(19) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(20) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(21) <= "0000000" & "00011" &"00000" &"010" & "00110" & "0100011";
-- mem(22) <= "0000000" & "00001" &"00000" &"010" & "00011" & "0100011";
-- mem(23) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(24) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(25) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(26) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(27) <= "0000000" & "00110" &"00000" &"010" & "01001" & "0000011";
-- mem(28) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(29) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(30) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(31) <= "0000000" & "00000" &"00000" &"000" & "00000" & "1100011";--beq r4,r5,-1
-- mem(32) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(33) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(34) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(35) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";



--mem(0) <= x"03000413";

--mem(1) <= x"04000793";
--mem(2) <= x"fef42623";

--mem(3) <= x"04400793";
--mem(4) <= x"fef42423";

--mem(5) <= x"04800793";
--mem(6) <= x"fef42223";

--mem(7) <= x"fe842783";
--mem(8) <= x"00a00713";
--mem(9) <= x"00e7a023";

--mem(10)<= x"fec42783";
--mem(11)<= x"00300713";
--mem(12)<= x"00e7a023";

--mem(13)<= x"fec42783";
--mem(14)<= x"00000033";
--mem(15)<= x"0007a703";
--mem(16)<= x"00000033";
--mem(17)<= x"fe842783";
--mem(18)<= x"00000033";
--mem(19)<= x"0007a783";
--mem(20)<= x"00000033";
--mem(21)<= x"00f70733";
--mem(22)<= x"fe442783";
--mem(23)<= x"00000033";
--mem(24)<= x"00e7a023";
--mem(25)<= x"0000006f";
--mem(26)<= x"0000006f";
--mem(27)<= x"0000006f";
--mem(28)<= x"0000006f";
--mem(29)<= x"0000006f";

    o_data <= mem(to_integer(unsigned(( i_addr(31 downto 2)))));
    o_valid<='1';
end behave;

--   10114:	01000793          	li	a5,16
--   10118:	fef42623          	sw	a5,-20(s0)
--   1011c:	01400793          	li	a5,20
--   10120:	fef42423          	sw	a5,-24(s0)
--   10124:	01800793          	li	a5,24
--   10128:	fef42223          	sw	a5,-28(s0)
--   1012c:	fe842783          	lw	a5,-24(s0)
--   10130:	00a00713          	li	a4,10
--   10134:	00e7a023          	sw	a4,0(a5)
--   10138:	fec42783          	lw	a5,-20(s0)
--   1013c:	00300713          	li	a4,3
--   10140:	00e7a023          	sw	a4,0(a5)
--   10144:	fec42783          	lw	a5,-20(s0)
--   10148:	0007a703          	lw	a4,0(a5)
--   1014c:	fe842783          	lw	a5,-24(s0)
--   10150:	0007a783          	lw	a5,0(a5)
--   10154:	00f70733          	add	a4,a4,a5
--   10158:	fe442783          	lw	a5,-28(s0)
--   1015c:	00e7a023          	sw	a4,0(a5)
--   10160:	0000006f          	j	10160 <main+0
