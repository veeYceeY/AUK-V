----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10.05.2020 11:12:15
-- Design Name: 
-- Module Name: pkg_sciv - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
package pkg_sciv is

constant LUI : std_logic_vector(7 downto 0)     := "00110111";
constant AUIPC : std_logic_vector(7 downto 0)   := "00010111";
constant JAL : std_logic_vector(7 downto 0)     := "01101111";
constant JALR : std_logic_vector(7 downto 0) := "0110011";
constant BEQ : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";
constant LUIPC : std_logic_vector(7 downto 0) := "00110111";

end package;