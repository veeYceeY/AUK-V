library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;


entity code_mem is
    port(
            i_en : in std_logic;
            i_addr : in std_logic_vector(31 downto 0);
            o_data : out std_logic_vector(31 downto 0);
            o_valid: out std_logic
    );

end code_mem;

architecture behave of code_mem is
type mem_type is array(63 downto 0) of std_logic_vector(31 downto 0);
signal mem : mem_type;

begin

--     --        
     
-- mem(0) <= x"00044" & "00100" & "0110111";--LUI r1,#00044000h
-- mem(1) <= x"00032" & "00101" & "0110111";--LUI r2,#00032000h
-- mem(2) <= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R1,12
-- mem(3) <= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R2,12
-- mem(4) <= "0000000" & "00101" &"00100" &"000" & "00011" & "0110011";--ADD r3,r1,r2
-- mem(5) <= x"0000a" & "00001" & "0110111";--LUI r1,#00044000h
-- mem(6) <= x"00003" & "00010" & "0110111";--LUI r2,#00032000h
-- mem(7) <= "0000000" & "01100" &"00001" &"101" & "00001" & "0010011";--srlI R1,12
-- mem(8) <= "0000000" & "01100" &"00010" &"101" & "00010" & "0010011";--srlI R2,12
-- mem(9) <= x"0000f" & "00100" & "0110111";--LUI r4,0x0000a000
-- mem(10)<= x"00002" & "00101" & "0110111";--LUI r5,0x00004000
-- mem(11)<= x"00001" & "00110" & "0110111";--LUI r6,0x00001000
-- mem(12)<= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R4,12
-- mem(13)<= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R5,12
-- mem(14) <="0000000" & "01100" &"00110" &"101" & "00110" & "0010011";--srlI R6,12
-- mem(15) <= "0100000" & "00110" &"00100" &"000" & "00100" & "0110011";--sub r4,r4,r6
-- mem(16) <= "1111111" & "00100" &"00101" &"100" & "11101" & "1100011";--blt r4,r5,-1
-- mem(17) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(18) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(19) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(20) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(21) <= "0000000" & "00011" &"00000" &"010" & "00110" & "0100011";
-- mem(22) <= "0000000" & "00001" &"00000" &"010" & "00011" & "0100011";
-- mem(23) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(24) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(25) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(26) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(27) <= "0000000" & "00110" &"00000" &"010" & "01001" & "0000011";
-- mem(28) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(29) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(30) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(31) <= "0000000" & "00000" &"00000" &"000" & "00000" & "1100011";--beq r4,r5,-1
-- mem(32) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(33) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(34) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(35) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";


mem(0) <= x"00812e23";
mem(1) <= x"02010413";
mem(2) <= x"00a00793";
mem(3) <= x"fef42623";
mem(4) <= x"03000793";
mem(5) <= x"fef42423";
mem(6) <= x"fe040793";
mem(7) <= x"fef42223";
mem(8) <= x"fe442783";
mem(9) <= x"00800713";
mem(10)<= x"00e7a023";
mem(11)<= x"0000006f";
mem(12)<= x"fe010113";
mem(13)<= x"fe010113";
mem(14)<= x"fe010113";
mem(15)<= x"fe010113";
mem(16)<= x"fe010113";

    o_data <= mem(to_integer(unsigned(( i_addr(31 downto 2)))));
    o_valid<='1';
end behave;


-- 10108:	fe010113          	addi	sp,sp,-32
--    1010c:	00812e23          	sw	s0,28(sp)
--    10110:	02010413          	addi	s0,sp,32
-- /home/veeyceey/eclipse-workspace/td/Debug/../src/main.cpp:26
--  // cout << "Hello RISC-V World!" << endl;
--   int gpio;
--   int *ptr;
--   int a,b,c;
--   b=10;
--    10114:	00a00793          	li	a5,10
--    10118:	fef42623          	sw	a5,-20(s0)
-- /home/veeyceey/eclipse-workspace/td/Debug/../src/main.cpp:27
--   a=48;
--    1011c:	03000793          	li	a5,48
--    10120:	fef42423          	sw	a5,-24(s0)
-- /home/veeyceey/eclipse-workspace/td/Debug/../src/main.cpp:29
--   //c=a*b;
--   ptr =&gpio;
--    10124:	fe040793          	addi	a5,s0,-32
--    10128:	fef42223          	sw	a5,-28(s0)
-- /home/veeyceey/eclipse-workspace/td/Debug/../src/main.cpp:30
--   *ptr=0x0008;
--    1012c:	fe442783          	lw	a5,-28(s0)
--    10130:	00800713          	li	a4,8
--    10134:	00e7a023          	sw	a4,0(a5)
-- /home/veeyceey/eclipse-workspace/td/Debug/../src/main.cpp:31 (discriminator 1)
--   while(1){}
--    10138:	0000006f          	j	10138 <main+0x30>


--    00812e23
--    02010413
--    00a00793
--    fef42623
--    03000793
--    fef42423
--    fe040793
--    fef42223
--    fe442783
--    00800713
--    00e7a023
--    0000006f




