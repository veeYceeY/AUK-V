library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;


entity code_mem is
    port(
            i_en : in std_logic;
            i_addr : in std_logic_vector(31 downto 0);
            o_data : out std_logic_vector(31 downto 0);
            o_valid: out std_logic
    );

end code_mem;

architecture behave of code_mem is
attribute rom_style : string;
type mem_type is array(511 downto 0) of std_logic_vector(31 downto 0);
signal mem : mem_type;
attribute rom_style of mem : signal is "block";

begin
--mem(0) <=x"03000413";
--mem(1) <=x"04000793";
--mem(2) <=x"FEF42623";
--mem(3) <=x"04400793";
--mem(4) <=x"FEF42423";
--mem(5) <=x"04800793";
--mem(6) <=x"FEF42223";
--mem(7) <=x"FE842783";
--mem(8) <=x"00A00713";
--mem(9) <=x"00E7A023";
--mem(10)<=x"FEC42783";
--mem(11)<=x"00400713";
--mem(12)<=x"00E7A023";
--mem(13)<=x"FEC42783";
--mem(14)<=x"0007A703";
--mem(15)<=x"FE842783";
--mem(16)<=x"0007A783";
--mem(17)<=x"00F70733";
--mem(18)<=x"FE442783";
--mem(19)<=x"00E7A023";
--mem(20)<=x"0000006F";

--working woith loops ---------
mem(54)<=x"03000413";--
mem(55)<=x"04000793";
mem(56)<=x"FEF42023";
mem(57)<=x"04400793";
mem(58)<=x"FCF42E23";
mem(59)<=x"04800793";
mem(60)<=x"FCF42C23";
mem(61)<=x"FE042783";
mem(62)<=x"00500713";
mem(63)<=x"00E7A023";
mem(64)<=x"FDC42783";
mem(65)<=x"00A00713";
mem(66)<=x"00E7A023";
mem(67)<=x"FE042783";
mem(68)<=x"0007A703";
mem(69)<=x"FDC42783";
mem(70)<=x"0007A783";
mem(71)<=x"00F70733";
mem(72)<=x"FD842783";
mem(73)<=x"00E7A023";
mem(74)<=x"000017B7";
mem(75)<=x"00178793";
mem(76)<=x"FCF42A23";
mem(77)<=x"FD442783";
mem(78)<=x"08600713";
mem(79)<=x"00E7A023";
mem(80)<=x"FE042623";
mem(81)<=x"FEC42703";
mem(82)<=x"0007A7B7";
mem(83)<=x"11F78793";
mem(84)<=x"00E7CA63";
mem(85)<=x"FEC42783";
mem(86)<=x"00178793";
mem(87)<=x"FEF42623";
mem(88)<=x"FE5FF06F";
mem(89)<=x"FD442783";
mem(90)<=x"04500713";
mem(91)<=x"00E7A023";
mem(92)<=x"FE042423";
mem(93)<=x"FE842703";
mem(94)<=x"0007A7B7";
mem(95)<=x"11F78793";
mem(96)<=x"00E7CA63";
mem(97)<=x"FE842783";
mem(98)<=x"00178793";
mem(99)<=x"FEF42423";
mem(100)<=x"FE5FF06F";
mem(101)<=x"FD442783";
mem(102)<=x"07600713";
mem(103)<=x"00E7A023";
mem(104)<=x"FE042223";
mem(105)<=x"FE442703";
mem(106)<=x"0007A7B7";
mem(107)<=x"11F78793";
mem(108)<=x"00E7CA63";
mem(109)<=x"FE442783";
mem(110)<=x"00178793";
mem(111)<=x"FEF42223";
mem(112)<=x"FE5FF06F";
mem(113)<=x"FD442783";
mem(114)<=x"0E300713";
mem(115)<=x"00E7A023";
mem(116)<=x"F71FF06F";





--mem(0) <=x"03000413";
--mem(1) <=x"FEF42423";--
--mem(2) <=x"04400793";
--mem(3) <=x"FEF42223";
--mem(4) <=x"04800793";
--mem(5) <=x"FEF42023";
--mem(6) <=x"FE442783";
--mem(7) <=x"00A00713";
--mem(8) <=x"00E7A023";
--mem(9) <=x"FE842783";
--mem(10)<=x"00400713";
--mem(11)<=x"00E7A023";
--mem(12)<=x"FE842783";
--mem(13)<=x"0007A703";
--mem(14)<=x"FE442783";
--mem(15)<=x"0007A783";
--mem(16)<=x"00F70733";
--mem(17)<=x"FE042783";
--mem(18)<=x"00E7A023";
--mem(19)<=x"04C00793";
--mem(20)<=x"FCF42E23";
--mem(21)<=x"FDC42783";
--mem(22)<=x"0007A023";
--mem(23)<=x"FE042623";
--mem(24)<=x"FE442783";
--mem(25)<=x"0007A783";
--mem(26)<=x"FEC42703";
--mem(27)<=x"02F75863";
--mem(28)<=x"FE842783";
--mem(29)<=x"0007A703";
--mem(30)<=x"FDC42783";
--mem(31)<=x"0007A783";
--mem(32)<=x"00F70733";
--mem(33)<=x"FDC42783";
--mem(34)<=x"00E7A023";
--mem(35)<=x"FEC42783";
--mem(36)<=x"00178793";
--mem(37)<=x"FEF42623";
--mem(38)<=x"FC9FF06F";
--mem(39)<=x"0000006F";-----


--mem(0)<=x"00000793";
--mem(1)<=x"00078863";
--mem(2)<=x"00010537";
--mem(3)<=x"46850513";
--mem(4)<=x"4400006F";
--mem(5)<=x"00008067";
--mem(6)<=x"00002197";
--mem(7)<=x"D7418193";
--mem(8)<=x"C3018513";
--mem(9)<=x"C4C18613";
--mem(10)<=x"40A60633";
--mem(11)<=x"00000593";
--mem(12)<=x"1C8000EF";
--mem(13)<=x"00000517";
--mem(14)<=x"41C50513";
--mem(15)<=x"00050863";
--mem(16)<=x"00000517";
--mem(17)<=x"3B450513";
--mem(18)<=x"408000EF";
--mem(19)<=x"110000EF";
--mem(20)<=x"00012503";
--mem(21)<=x"00410593";
--mem(22)<=x"00000613";
--mem(23)<=x"074000EF";
--mem(24)<=x"0CC0006F";
--mem(25)<=x"C301C703";
--mem(26)<=x"04071263";
--mem(27)<=x"FF010113";
--mem(28)<=x"00812423";
--mem(29)<=x"00078413";
--mem(30)<=x"00112623";
--mem(31)<=x"00000793";
--mem(32)<=x"00078A63";
--mem(33)<=x"00011537";
--mem(34)<=x"5BC50513";
--mem(35)<=x"00000097";
--mem(36)<=x"000000E7";
--mem(37)<=x"00100793";
--mem(38)<=x"00C12083";
--mem(39)<=x"C2F18823";
--mem(40)<=x"00812403";
--mem(41)<=x"01010113";
--mem(42)<=x"00008067";
--mem(43)<=x"00008067";
--mem(44)<=x"00000793";
--mem(45)<=x"00078C63";
--mem(46)<=x"00011537";
--mem(47)<=x"C3418593";
--mem(48)<=x"5BC50513";
--mem(49)<=x"00000317";
--mem(50)<=x"00000067";
--mem(51)<=x"00008067";
--mem(52)<=x"FE010113";
--mem(53)<=x"00812E23";
--mem(54)<=x"02010413";
--mem(55)<=x"04000793";
--mem(56)<=x"FEF42623";
--mem(57)<=x"04400793";
--mem(58)<=x"FEF42423";
--mem(59)<=x"04800793";
--mem(60)<=x"FEF42223";
--mem(61)<=x"FE842783";
--mem(62)<=x"00A00713";
--mem(63)<=x"00E7A023";
--mem(64)<=x"FEC42783";
--mem(65)<=x"00400713";
--mem(66)<=x"00E7A023";
--mem(67)<=x"FEC42783";
--mem(68)<=x"0007A703";
--mem(69)<=x"FE842783";
--mem(70)<=x"0007A783";
--mem(71)<=x"00F70733";
--mem(72)<=x"FE442783";
--mem(73)<=x"00E7A023";
--mem(74)<=x"0000006F";
--mem(75)<=x"FF010113";
--mem(76)<=x"00000593";
--mem(77)<=x"00812423";
--mem(78)<=x"00112623";
--mem(79)<=x"00050413";
--mem(80)<=x"194000EF";
--mem(81)<=x"C281A503";
--mem(82)<=x"03C52783";
--mem(83)<=x"00078463";
--mem(84)<=x"000780E7";
--mem(85)<=x"00040513";
--mem(86)<=x"3A4000EF";
--mem(87)<=x"FF010113";
--mem(88)<=x"00812423";
--mem(89)<=x"01212023";
--mem(90)<=x"00011437";
--mem(91)<=x"00011937";
--mem(92)<=x"5F040793";
--mem(93)<=x"5F090913";
--mem(94)<=x"40F90933";
--mem(95)<=x"00112623";
--mem(96)<=x"00912223";
--mem(97)<=x"40295913";
--mem(98)<=x"02090063";
--mem(99)<=x"5F040413";
--mem(100)<=x"00000493";
--mem(101)<=x"00042783";
--mem(102)<=x"00148493";
--mem(103)<=x"00440413";
--mem(104)<=x"000780E7";
--mem(105)<=x"FE9918E3";
--mem(106)<=x"00011437";
--mem(107)<=x"00011937";
--mem(108)<=x"5F040793";
--mem(109)<=x"5F890913";
--mem(110)<=x"40F90933";
--mem(111)<=x"40295913";
--mem(112)<=x"02090063";
--mem(113)<=x"5F040413";
--mem(114)<=x"00000493";
--mem(115)<=x"00042783";
--mem(116)<=x"00148493";
--mem(117)<=x"00440413";
--mem(118)<=x"000780E7";
--mem(119)<=x"FE9918E3";
--mem(120)<=x"00C12083";
--mem(121)<=x"00812403";
--mem(122)<=x"00412483";
--mem(123)<=x"00012903";
--mem(124)<=x"01010113";
--mem(125)<=x"00008067";
--mem(126)<=x"00F00313";
--mem(127)<=x"00050713";
--mem(128)<=x"02C37E63";
--mem(129)<=x"00F77793";
--mem(130)<=x"0A079063";
--mem(131)<=x"08059263";
--mem(132)<=x"FF067693";
--mem(133)<=x"00F67613";
--mem(134)<=x"00E686B3";
--mem(135)<=x"00B72023";
--mem(136)<=x"00B72223";
--mem(137)<=x"00B72423";
--mem(138)<=x"00B72623";
--mem(139)<=x"01070713";
--mem(140)<=x"FED766E3";
--mem(141)<=x"00061463";
--mem(142)<=x"00008067";
--mem(143)<=x"40C306B3";
--mem(144)<=x"00269693";
--mem(145)<=x"00000297";
--mem(146)<=x"005686B3";
--mem(147)<=x"00C68067";
--mem(148)<=x"00B70723";
--mem(149)<=x"00B706A3";
--mem(150)<=x"00B70623";
--mem(151)<=x"00B705A3";
--mem(152)<=x"00B70523";
--mem(153)<=x"00B704A3";
--mem(154)<=x"00B70423";
--mem(155)<=x"00B703A3";
--mem(156)<=x"00B70323";
--mem(157)<=x"00B702A3";
--mem(158)<=x"00B70223";
--mem(159)<=x"00B701A3";
--mem(160)<=x"00B70123";
--mem(161)<=x"00B700A3";
--mem(162)<=x"00B70023";
--mem(163)<=x"00008067";
--mem(164)<=x"0FF5F593";
--mem(165)<=x"00859693";
--mem(166)<=x"00D5E5B3";
--mem(167)<=x"01059693";
--mem(168)<=x"00D5E5B3";
--mem(169)<=x"F6DFF06F";
--mem(170)<=x"00279693";
--mem(171)<=x"00000297";
--mem(172)<=x"005686B3";
--mem(173)<=x"00008293";
--mem(174)<=x"FA0680E7";
--mem(175)<=x"00028093";
--mem(176)<=x"FF078793";
--mem(177)<=x"40F70733";
--mem(178)<=x"00F60633";
--mem(179)<=x"F6C378E3";
--mem(180)<=x"F3DFF06F";
--mem(181)<=x"FD010113";
--mem(182)<=x"01412C23";
--mem(183)<=x"C281AA03";
--mem(184)<=x"03212023";
--mem(185)<=x"02112623";
--mem(186)<=x"148A2903";
--mem(187)<=x"02812423";
--mem(188)<=x"02912223";
--mem(189)<=x"01312E23";
--mem(190)<=x"01512A23";
--mem(191)<=x"01612823";
--mem(192)<=x"01712623";
--mem(193)<=x"01812423";
--mem(194)<=x"04090063";
--mem(195)<=x"00050B13";
--mem(196)<=x"00058B93";
--mem(197)<=x"00100A93";
--mem(198)<=x"FFF00993";
--mem(199)<=x"00492483";
--mem(200)<=x"FFF48413";
--mem(201)<=x"02044263";
--mem(202)<=x"00249493";
--mem(203)<=x"009904B3";
--mem(204)<=x"040B8463";
--mem(205)<=x"1044A783";
--mem(206)<=x"05778063";
--mem(207)<=x"FFF40413";
--mem(208)<=x"FFC48493";
--mem(209)<=x"FF3416E3";
--mem(210)<=x"02C12083";
--mem(211)<=x"02812403";
--mem(212)<=x"02412483";
--mem(213)<=x"02012903";
--mem(214)<=x"01C12983";
--mem(215)<=x"01812A03";
--mem(216)<=x"01412A83";
--mem(217)<=x"01012B03";
--mem(218)<=x"00C12B83";
--mem(219)<=x"00812C03";
--mem(220)<=x"03010113";
--mem(221)<=x"00008067";
--mem(222)<=x"00492783";
--mem(223)<=x"0044A683";
--mem(224)<=x"FFF78793";
--mem(225)<=x"04878E63";
--mem(226)<=x"0004A223";
--mem(227)<=x"FA0688E3";
--mem(228)<=x"18892783";
--mem(229)<=x"008A9733";
--mem(230)<=x"00492C03";
--mem(231)<=x"00F777B3";
--mem(232)<=x"02079263";
--mem(233)<=x"000680E7";
--mem(234)<=x"00492703";
--mem(235)<=x"148A2783";
--mem(236)<=x"01871463";
--mem(237)<=x"F92784E3";
--mem(238)<=x"F80788E3";
--mem(239)<=x"00078913";
--mem(240)<=x"F5DFF06F";
--mem(241)<=x"18C92783";
--mem(242)<=x"0844A583";
--mem(243)<=x"00F77733";
--mem(244)<=x"00071C63";
--mem(245)<=x"000B0513";
--mem(246)<=x"000680E7";
--mem(247)<=x"FCDFF06F";
--mem(248)<=x"00892223";
--mem(249)<=x"FA9FF06F";
--mem(250)<=x"00058513";
--mem(251)<=x"000680E7";
--mem(252)<=x"FB9FF06F";
--mem(253)<=x"FF010113";
--mem(254)<=x"00812423";
--mem(255)<=x"000117B7";
--mem(256)<=x"00011437";
--mem(257)<=x"5F840413";
--mem(258)<=x"5FC78793";
--mem(259)<=x"408787B3";
--mem(260)<=x"00912223";
--mem(261)<=x"00112623";
--mem(262)<=x"4027D493";
--mem(263)<=x"02048063";
--mem(264)<=x"FFC78793";
--mem(265)<=x"00878433";
--mem(266)<=x"00042783";
--mem(267)<=x"FFF48493";
--mem(268)<=x"FFC40413";
--mem(269)<=x"000780E7";
--mem(270)<=x"FE0498E3";
--mem(271)<=x"00C12083";
--mem(272)<=x"00812403";
--mem(273)<=x"00412483";
--mem(274)<=x"01010113";
--mem(275)<=x"00008067";
--mem(276)<=x"00050593";
--mem(277)<=x"00000693";
--mem(278)<=x"00000613";
--mem(279)<=x"00000513";
--mem(280)<=x"0040006F";
--mem(281)<=x"C281A703";
--mem(282)<=x"14872783";
--mem(283)<=x"04078C63";
--mem(284)<=x"0047A703";
--mem(285)<=x"01F00813";
--mem(286)<=x"06E84E63";
--mem(287)<=x"00271813";
--mem(288)<=x"02050663";
--mem(289)<=x"01078333";
--mem(290)<=x"08C32423";
--mem(291)<=x"1887A883";
--mem(292)<=x"00100613";
--mem(293)<=x"00E61633";
--mem(294)<=x"00C8E8B3";
--mem(295)<=x"1917A423";
--mem(296)<=x"10D32423";
--mem(297)<=x"00200693";
--mem(298)<=x"02D50463";
--mem(299)<=x"00170713";
--mem(300)<=x"00E7A223";
--mem(301)<=x"010787B3";
--mem(302)<=x"00B7A423";
--mem(303)<=x"00000513";
--mem(304)<=x"00008067";
--mem(305)<=x"14C70793";
--mem(306)<=x"14F72423";
--mem(307)<=x"FA5FF06F";
--mem(308)<=x"18C7A683";
--mem(309)<=x"00170713";
--mem(310)<=x"00E7A223";
--mem(311)<=x"00C6E633";
--mem(312)<=x"18C7A623";
--mem(313)<=x"010787B3";
--mem(314)<=x"00B7A423";
--mem(315)<=x"00000513";
--mem(316)<=x"00008067";
--mem(317)<=x"FFF00513";
--mem(318)<=x"00008067";
--mem(319)<=x"00000593";
--mem(320)<=x"00000613";
--mem(321)<=x"00000693";
--mem(322)<=x"00000713";
--mem(323)<=x"00000793";
--mem(324)<=x"05D00893";
--mem(325)<=x"00000073";
--mem(326)<=x"00054463";
--mem(327)<=x"0000006F";
--mem(328)<=x"FF010113";
--mem(329)<=x"00812423";
--mem(330)<=x"00050413";
--mem(331)<=x"00112623";
--mem(332)<=x"40800433";
--mem(333)<=x"00C000EF";
--mem(334)<=x"00852023";
--mem(335)<=x"0000006F";
--mem(336)<=x"C2C1A503";
--mem(337)<=x"00008067";
--mem(338)<=x"00000010";
--mem(339)<=x"00000000";
--mem(340)<=x"00527A03";
--mem(341)<=x"01017C01";
--mem(342)<=x"00020D1B";
--mem(343)<=x"00000018";
--mem(344)<=x"00000018";
--mem(345)<=x"FFFFEB6C";
--mem(346)<=x"0000005C";
--mem(347)<=x"200E4400";
--mem(348)<=x"44018844";
--mem(349)<=x"0000080C";
--mem(350)<=x"00000000";
--mem(351)<=x"00010074";
--mem(352)<=x"00010124";
--mem(353)<=x"000100D8";
--mem(354)<=x"00000000";
--mem(355)<=x"000118EC";
--mem(356)<=x"00011954";
--mem(357)<=x"000119BC";
--mem(358)<=x"00000000";
--mem(359)<=x"00000000";
--mem(360)<=x"00000000";
--mem(361)<=x"00000000";
--mem(362)<=x"00000000";
--mem(363)<=x"00000000";
--mem(364)<=x"00000000";
--mem(365)<=x"00000000";
--mem(366)<=x"00000000";
--mem(367)<=x"00000000";
--mem(368)<=x"00000000";
--mem(369)<=x"00000000";
--mem(370)<=x"00000000";
--mem(371)<=x"00000000";
--mem(372)<=x"00000000";
--mem(373)<=x"00000000";
--mem(374)<=x"00000000";
--mem(375)<=x"00000000";
--mem(376)<=x"00000000";
--mem(377)<=x"00000000";
--mem(378)<=x"00000000";
--mem(379)<=x"00000000";
--mem(380)<=x"00000000";
--mem(381)<=x"00000000";
--mem(382)<=x"00000000";
--mem(383)<=x"00000000";
--mem(384)<=x"00000000";
--mem(385)<=x"00000000";
--mem(386)<=x"00000000";
--mem(387)<=x"00000000";
--mem(388)<=x"00000000";
--mem(389)<=x"00000000";
--mem(390)<=x"00000000";
--mem(391)<=x"00000000";
--mem(392)<=x"00000000";
--mem(393)<=x"00000000";
--mem(394)<=x"00000000";
--mem(395)<=x"00000000";
--mem(396)<=x"00000001";
--mem(397)<=x"00000000";
--mem(398)<=x"ABCD330E";
--mem(399)<=x"E66D1234";
--mem(400)<=x"0005DEEC";
--mem(401)<=x"0000000B";
--mem(402)<=x"00000000";
--mem(403)<=x"00000000";
--mem(404)<=x"00000000";
--mem(405)<=x"00000000";
--mem(406)<=x"00000000";
--mem(407)<=x"00000000";
--mem(408)<=x"00000000";
--mem(409)<=x"00000000";
--mem(410)<=x"00000000";
--mem(411)<=x"00000000";
--mem(412)<=x"00000000";
--mem(413)<=x"00000000";
--mem(414)<=x"00000000";
--mem(415)<=x"00000000";
--mem(416)<=x"00000000";
--mem(417)<=x"00000000";
--mem(418)<=x"00000000";
--mem(419)<=x"00000000";
--mem(420)<=x"00000000";
--mem(421)<=x"00000000";
--mem(422)<=x"00000000";
--mem(423)<=x"00000000";
--mem(424)<=x"00000000";
--mem(425)<=x"00000000";
--mem(426)<=x"00000000";
--mem(427)<=x"00000000";
--mem(428)<=x"00000000";
--mem(429)<=x"00000000";
--mem(430)<=x"00000000";
--mem(431)<=x"00000000";
--mem(432)<=x"00000000";
--mem(433)<=x"00000000";
--mem(434)<=x"00000000";
--mem(435)<=x"00000000";
--mem(436)<=x"00000000";
--mem(437)<=x"00000000";
--mem(438)<=x"00000000";
--mem(439)<=x"00000000";
--mem(440)<=x"00000000";
--mem(441)<=x"00000000";
--mem(442)<=x"00000000";
--mem(443)<=x"00000000";
--mem(444)<=x"00000000";
--mem(445)<=x"00000000";
--mem(446)<=x"00000000";
--mem(447)<=x"00000000";
--mem(448)<=x"00000000";
--mem(449)<=x"00000000";
--mem(450)<=x"00000000";
--mem(451)<=x"00000000";
--mem(452)<=x"00000000";
--mem(453)<=x"00000000";
--mem(454)<=x"00000000";
--mem(455)<=x"00000000";
--mem(456)<=x"00000000";
--mem(457)<=x"00000000";
--mem(458)<=x"00000000";
--mem(459)<=x"00000000";
--mem(460)<=x"00000000";
--mem(461)<=x"00000000";
--mem(462)<=x"00000000";
--mem(463)<=x"00000000";
--mem(464)<=x"00000000";
--mem(465)<=x"00000000";
--mem(466)<=x"00000000";
--mem(467)<=x"00000000";
--mem(468)<=x"00000000";
--mem(469)<=x"00000000";
--mem(470)<=x"00000000";
--mem(471)<=x"00000000";
--mem(472)<=x"00000000";
--mem(473)<=x"00000000";
--mem(474)<=x"00000000";
--mem(475)<=x"00000000";
--mem(476)<=x"00000000";
--mem(477)<=x"00000000";
--mem(478)<=x"00000000";
--mem(479)<=x"00000000";
--mem(480)<=x"00000000";
--mem(481)<=x"00000000";
--mem(482)<=x"00000000";
--mem(483)<=x"00000000";
--mem(484)<=x"00000000";
--mem(485)<=x"00000000";
--mem(486)<=x"00000000";
--mem(487)<=x"00000000";
--mem(488)<=x"00000000";
--mem(489)<=x"00000000";
--mem(490)<=x"00000000";
--mem(491)<=x"00000000";
--mem(492)<=x"00000000";
--mem(493)<=x"00000000";
--mem(494)<=x"00000000";
--mem(495)<=x"00000000";
--mem(496)<=x"00000000";
--mem(497)<=x"00000000";
--mem(498)<=x"00000000";
--mem(499)<=x"00000000";
--mem(500)<=x"00000000";
--mem(501)<=x"00000000";
--mem(502)<=x"00000000";
--mem(503)<=x"00000000";
--mem(504)<=x"00000000";
--mem(505)<=x"00000000";
--mem(506)<=x"00000000";
--mem(507)<=x"00000000";
--mem(508)<=x"00000000";
--mem(509)<=x"00000000";
--mem(510)<=x"00000000";
--mem(511)<=x"00000000";
--mem(512)<=x"00000000";
--mem(513)<=x"00000000";
--mem(514)<=x"00000000";
--mem(515)<=x"00000000";
--mem(516)<=x"00000000";
--mem(517)<=x"00000000";
--mem(518)<=x"00000000";
--mem(519)<=x"00000000";
--mem(520)<=x"00000000";
--mem(521)<=x"00000000";
--mem(522)<=x"00000000";
--mem(523)<=x"00000000";
--mem(524)<=x"00000000";
--mem(525)<=x"00000000";
--mem(526)<=x"00000000";
--mem(527)<=x"00000000";
--mem(528)<=x"00000000";
--mem(529)<=x"00000000";
--mem(530)<=x"00000000";
--mem(531)<=x"00000000";
--mem(532)<=x"00000000";
--mem(533)<=x"00000000";
--mem(534)<=x"00000000";
--mem(535)<=x"00000000";
--mem(536)<=x"00000000";
--mem(537)<=x"00000000";
--mem(538)<=x"00000000";
--mem(539)<=x"00000000";
--mem(540)<=x"00000000";
--mem(541)<=x"00000000";
--mem(542)<=x"00000000";
--mem(543)<=x"00000000";
--mem(544)<=x"00000000";
--mem(545)<=x"00000000";
--mem(546)<=x"00000000";
--mem(547)<=x"00000000";
--mem(548)<=x"00000000";
--mem(549)<=x"00000000";
--mem(550)<=x"00000000";
--mem(551)<=x"00000000";
--mem(552)<=x"00000000";
--mem(553)<=x"00000000";
--mem(554)<=x"00000000";
--mem(555)<=x"00000000";
--mem(556)<=x"00000000";
--mem(557)<=x"00000000";
--mem(558)<=x"00000000";
--mem(559)<=x"00000000";
--mem(560)<=x"00000000";
--mem(561)<=x"00000000";
--mem(562)<=x"00000000";
--mem(563)<=x"00000000";
--mem(564)<=x"00000000";
--mem(565)<=x"00000000";
--mem(566)<=x"00000000";
--mem(567)<=x"00000000";
--mem(568)<=x"00000000";
--mem(569)<=x"00000000";
--mem(570)<=x"00000000";
--mem(571)<=x"00000000";
--mem(572)<=x"00000000";
--mem(573)<=x"00000000";
--mem(574)<=x"00000000";
--mem(575)<=x"00000000";
--mem(576)<=x"00000000";
--mem(577)<=x"00000000";
--mem(578)<=x"00000000";
--mem(579)<=x"00000000";
--mem(580)<=x"00000000";
--mem(581)<=x"00000000";
--mem(582)<=x"00000000";
--mem(583)<=x"00000000";
--mem(584)<=x"00000000";
--mem(585)<=x"00000000";
--mem(586)<=x"00000000";
--mem(587)<=x"00000000";
--mem(588)<=x"00000000";
--mem(589)<=x"00000000";
--mem(590)<=x"00000000";
--mem(591)<=x"00000000";
--mem(592)<=x"00000000";
--mem(593)<=x"00000000";
--mem(594)<=x"00000000";
--mem(595)<=x"00000000";
--mem(596)<=x"00000000";
--mem(597)<=x"00000000";
--mem(598)<=x"00000000";
--mem(599)<=x"00000000";
--mem(600)<=x"00000000";
--mem(601)<=x"00000000";
--mem(602)<=x"00000000";
--mem(603)<=x"00000000";
--mem(604)<=x"00000000";
--mem(605)<=x"00000000";
--mem(606)<=x"00000000";
--mem(607)<=x"00000000";
--mem(608)<=x"00000000";
--mem(609)<=x"00000000";
--mem(610)<=x"00000000";
--mem(611)<=x"00000000";
--mem(612)<=x"00000000";
--mem(613)<=x"00000000";
--mem(614)<=x"00000000";
--mem(615)<=x"00000000";
--mem(616)<=x"00000000";
--mem(617)<=x"00000000";
--mem(618)<=x"00000000";
--mem(619)<=x"00000000";
--mem(620)<=x"00011600";
--mem(621)<=x"00011600";

--     --        
     
-- mem(0) <= x"00044" & "00100" & "0110111";--LUI r1,#00044000h
-- mem(1) <= x"00032" & "00101" & "0110111";--LUI r2,#00032000h
-- mem(2) <= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R1,12
-- mem(3) <= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R2,12
-- mem(4) <= "0000000" & "00101" &"00100" &"000" & "00011" & "0110011";--ADD r3,r1,r2
-- mem(5) <= x"0000a" & "00001" & "0110111";--LUI r1,#00044000h
-- mem(6) <= x"00003" & "00010" & "0110111";--LUI r2,#00032000h
-- mem(7) <= "0000000" & "01100" &"00001" &"101" & "00001" & "0010011";--srlI R1,12
-- mem(8) <= "0000000" & "01100" &"00010" &"101" & "00010" & "0010011";--srlI R2,12
-- mem(9) <= x"0000f" & "00100" & "0110111";--LUI r4,0x0000a000
-- mem(10)<= x"00002" & "00101" & "0110111";--LUI r5,0x00004000
-- mem(11)<= x"00001" & "00110" & "0110111";--LUI r6,0x00001000
-- mem(12)<= "0000000" & "01100" &"00100" &"101" & "00100" & "0010011";--srlI R4,12
-- mem(13)<= "0000000" & "01100" &"00101" &"101" & "00101" & "0010011";--srlI R5,12
-- mem(14) <="0000000" & "01100" &"00110" &"101" & "00110" & "0010011";--srlI R6,12
-- mem(15) <= "0100000" & "00110" &"00100" &"000" & "00100" & "0110011";--sub r4,r4,r6
-- mem(16) <= "1111111" & "00100" &"00101" &"100" & "11101" & "1100011";--blt r4,r5,-1
-- mem(17) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(18) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(19) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(20) <= "0000000" & "10000" &"10000" &"000" & "00000" & "0110011";
-- mem(21) <= "0000000" & "00011" &"00000" &"010" & "00110" & "0100011";
-- mem(22) <= "0000000" & "00001" &"00000" &"010" & "00011" & "0100011";
-- mem(23) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(24) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(25) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(26) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(27) <= "0000000" & "00110" &"00000" &"010" & "01001" & "0000011";
-- mem(28) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(29) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(30) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(31) <= "0000000" & "00000" &"00000" &"000" & "00000" & "1100011";--beq r4,r5,-1
-- mem(32) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(33) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(34) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";
-- mem(35) <= "0000000" & "00000" &"00000" &"000" & "00000" & "0110011";



--mem(0) <= x"03000413";

--mem(1) <= x"04000793";
--mem(2) <= x"fef42623";

--mem(3) <= x"04400793";
--mem(4) <= x"fef42423";

--mem(5) <= x"04800793";
--mem(6) <= x"fef42223";

--mem(7) <= x"fe842783";
--mem(8) <= x"00a00713";
--mem(9) <= x"00e7a023";

--mem(10)<= x"fec42783";
--mem(11)<= x"00300713";
--mem(12)<= x"00e7a023";

--mem(13)<= x"fec42783";
--mem(14)<= x"00000033";
--mem(15)<= x"0007a703";
--mem(16)<= x"00000033";
--mem(17)<= x"fe842783";
--mem(18)<= x"00000033";
--mem(19)<= x"0007a783";
--mem(20)<= x"00000033";
--mem(21)<= x"00f70733";
--mem(22)<= x"fe442783";
--mem(23)<= x"00000033";
--mem(24)<= x"00e7a023";
--mem(25)<= x"0000006f";
--mem(26)<= x"0000006f";
--mem(27)<= x"0000006f";
--mem(28)<= x"0000006f";
--mem(29)<= x"0000006f";

    o_data <= mem(to_integer(unsigned(( i_addr(31 downto 2)))));
    o_valid<='1';
end behave;

--   10114:	01000793          	li	a5,16
--   10118:	fef42623          	sw	a5,-20(s0)
--   1011c:	01400793          	li	a5,20
--   10120:	fef42423          	sw	a5,-24(s0)
--   10124:	01800793          	li	a5,24
--   10128:	fef42223          	sw	a5,-28(s0)
--   1012c:	fe842783          	lw	a5,-24(s0)
--   10130:	00a00713          	li	a4,10
--   10134:	00e7a023          	sw	a4,0(a5)
--   10138:	fec42783          	lw	a5,-20(s0)
--   1013c:	00300713          	li	a4,3
--   10140:	00e7a023          	sw	a4,0(a5)
--   10144:	fec42783          	lw	a5,-20(s0)
--   10148:	0007a703          	lw	a4,0(a5)
--   1014c:	fe842783          	lw	a5,-24(s0)
--   10150:	0007a783          	lw	a5,0(a5)
--   10154:	00f70733          	add	a4,a4,a5
--   10158:	fe442783          	lw	a5,-28(s0)
--   1015c:	00e7a023          	sw	a4,0(a5)
--   10160:	0000006f          	j	10160 <main+0
